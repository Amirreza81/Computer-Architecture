library verilog;
use verilog.vl_types.all;
entity AluC_Control_vlg_vec_tst is
end AluC_Control_vlg_vec_tst;
